LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE KSPackage IS

COMPONENT Adder IS
	PORT (
		A,B : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		Cin : IN  STD_LOGIC;
		Cout: OUT STD_LOGIC;
		Sum : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT RolComponent IS
	PORT (
		N      : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		OP     : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		RESULT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT ModulusAddition IS
	PORT (
		OpA, OpB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		Result: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT DeltaConstants IS
	PORT (
		ADDR : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
		DATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT RoundConstants IS
  PORT (
		ADDR : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		DATA : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT Mux2to1 IS
	PORT (
		A: IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		B: IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		S: IN  STD_LOGIC;
		C: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;


COMPONENT RAMMemory IS
	PORT (
		CLK		: IN  STD_LOGIC;
		ADDR 		: IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		WD			: IN  STD_LOGIC;
		DATA_IN	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_OUT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	 );
END COMPONENT;

COMPONENT BufferT IS
  PORT (
		CLK : IN  STD_LOGIC;
		WD	 : IN  STD_LOGIC;
		DATA_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATA_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	 );
END COMPONENT;

END KSPackage;

	
PACKAGE BODY KSPackage IS


 
END KSPackage;
