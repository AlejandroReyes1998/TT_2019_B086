LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_BIT.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Mux2to1 IS

	GENERIC (
		N : INTEGER := 32
	);
	PORT (
		A: IN  STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		B: IN  STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		S: IN  STD_LOGIC;
		C: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
 
END Mux2to1;

ARCHITECTURE MuxArchitecture OF Mux2to1 IS

BEGIN

	C <= A when S else B;
	
END MuxArchitecture;