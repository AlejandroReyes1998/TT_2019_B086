LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL;

ENTITY ROLComponent IS
	
	PORT (
		N      : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		OP     : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		RESULT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
 
END ROLComponent;

ARCHITECTURE ROLArchitecture OF ROLComponent IS

BEGIN

  RESULT <= STD_LOGIC_VECTOR(UNSIGNED(OP) ROL TO_INTEGER(UNSIGNED(N)));
	
END ROLArchitecture;