LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.MATH_REAL.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;


ENTITY DeltaConstants IS

  PORT (
	 ADDR 							: IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
	 DATA								: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	 );
	 
END DeltaConstants;
 
ARCHITECTURE DCArchitecture OF DeltaConstants IS

TYPE ROM_MEMORY IS ARRAY (0 to 7) OF STD_LOGIC_VECTOR (31 downto 0);

SIGNAL ROM : ROM_MEMORY := ("11000011111011111110100111011011",
									 "01000100011000100110101100000010",
									 "01111001111000100111110010001010",
									 "01111000110111110011000011101100",
									 "01110001010111101010010010011110",
									 "11000111100001011101101000001010",
									 "11100000010011101111001000101010",
									 "11100101110001000000100101010111");
									 
BEGIN

	DATA <= ROM(CONV_INTEGER(ADDR));

END DCARCHITECTURE;
